interface cuboid_inp_intf (input clk);

  logic [16-1:0] in_data;
  logic          in_valid;
  logic          in_start;

endinterface
