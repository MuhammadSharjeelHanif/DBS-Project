 interface cuboid_out_intf (input clk);

  logic  [32-1:0]  out_data;
  logic            out_start;
  logic            out_valid;

endinterface