module test(sum,a,b);
	input a,b;
	output sum;

	or o1(sum, a,b);

endmodule


