package complex_pkg;
 `include "uvm_macros.svh"
  import uvm_pkg::*;
	
  //configs
  `include "complex_config.sv"
  `include "common_config.sv"
  // Sequence Item
  `include "complexnum.sv"
  // Drivers
  `include "inp_driver.sv"
  // Monitor
  `include "inp_monitor.sv"
  `include "out_monitor.sv"
  // Agents 
  `include "inp_agent.sv"
  `include "out_agent.sv"
  // Scoreboard
  `include "scoreboard.sv"
  // Sequences
  `include "complex_sequence.sv"
  `include "inp_sequence.sv"
  // Enironment 
  `include "env.sv"
  // Tests
  `include "complex_base_test.sv"
  `include "../test/new_test/test.sv"
endpackage 